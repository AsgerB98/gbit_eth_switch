library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use std.textio.all;
use IEEE.std_logic_textio.all;


entity ram is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        
    );
end entity;